
// `define BFU_USE_KARATSUBER
// `define TFG_USE_KARATSUBER
// `define TFG_NO_USE_DSP
// `define NO_DSP_NUM 0
`define BARRET_BYPASS